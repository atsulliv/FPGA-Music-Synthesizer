// How to use:					
// 1. Edit the songs on the Enter Song sheet.					
// 2. Select this whole worksheet, copy it, and paste it into a new file.					
// 3. Save the file as song_rom.v.					
					
module song_rom (					
	input clk,				
	input [8:0] addr,				
	output reg [15:0] dout				
);					
					
	wire [15:0] memory [511:0];				
					
	always @(posedge clk)				
		dout = memory[addr];			
					
	assign memory[	  0	] =	{1'd0, 6'd48, 6'd12, 3'd0};	// Note: 4G#Ab
	assign memory[	  1	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	  2	] =	{1'd0, 6'd52, 6'd12, 3'd0};	// Note: 5C
	assign memory[	  3	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	  4	] =	{1'd0, 6'd47, 6'd12, 3'd0};	// Note: 4G
	assign memory[	  5	] =	{1'd0, 6'd40, 6'd24, 3'd0};	// Note: 3G#Ab
	assign memory[	  6	] =	{1'd0, 6'd36, 6'd24, 3'd0};	// Note: 4C
	assign memory[	  7	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	  8	] =	{1'd0, 6'd48, 6'd12, 3'd0};	// Note: 4G#Ab
	assign memory[	  9	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 10	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	 11	] =	{1'd0, 6'd33, 6'd24, 3'd0};	// Note: 3F
	assign memory[	 12	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 13	] =	{1'd0, 6'd47, 6'd12, 3'd0};	// Note: 4G
	assign memory[	 14	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 15	] =	{1'd0, 6'd43, 6'd12, 3'd0};	// Note: 4D#Eb
	assign memory[	 16	] =	{1'd0, 6'd40, 6'd24, 3'd0};	// Note: 4C
	assign memory[	 17	] =	{1'd0, 6'd36, 6'd24, 3'd0};	// Note: 3G#Ab
	assign memory[	 18	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 19	] =	{1'd0, 6'd42, 6'd12, 3'd0};	// Note: 4D
	assign memory[	 20	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 21	] =	{1'd0, 6'd39, 6'd24, 3'd0};	// Note: 4B
	assign memory[	 22	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 23	] =	{1'd0, 6'd45, 6'd24, 3'd0};	// Note: 4F
	assign memory[	 24	] =	{1'd0, 6'd42, 6'd24, 3'd0};	// Note: 4D
	assign memory[	 25	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 26	] =	{1'd0, 6'd39, 6'd24, 3'd0};	// Note: 4B
	assign memory[	 27	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 28	] =	{1'd0, 6'd45, 6'd24, 3'd0};	// Note: 4F
	assign memory[	 29	] =	{1'd0, 6'd41, 6'd24, 3'd0};	// Note: 4C#Db
	assign memory[	 30	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 31	] =	{1'd0, 6'd36, 6'd24, 3'd0};	// Note: 3G#Ab
	assign memory[	 32	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 33	] =	{1'd0, 6'd33, 6'd24, 3'd0};	// Note: 3F
	assign memory[	 34	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 35	] =	{1'd0, 6'd52, 6'd12, 3'd0};	// Note: 5C
	assign memory[	 36	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 37	] =	{1'd0, 6'd46, 6'd24, 3'd0};	// Note: 4F#Gb
	assign memory[	 38	] =	{1'd0, 6'd40, 6'd24, 3'd0};	// Note: 4C
	assign memory[	 39	] =	{1'd0, 6'd36, 6'd24, 3'd0};	// Note: 3G#Ab
	assign memory[	 40	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 41	] =	{1'd0, 6'd48, 6'd12, 3'd0};	// Note: 4G#Ab
	assign memory[	 42	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 43	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	 44	] =	{1'd0, 6'd33, 6'd24, 3'd0};	// Note: 3F
	assign memory[	 45	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 46	] =	{1'd0, 6'd47, 6'd12, 3'd0};	// Note: 4G
	assign memory[	 47	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 48	] =	{1'd0, 6'd48, 6'd12, 3'd0};	// Note: 4G#Ab
	assign memory[	 49	] =	{1'd0, 6'd40, 6'd24, 3'd0};	// Note: 4C
	assign memory[	 50	] =	{1'd0, 6'd36, 6'd24, 3'd0};	// Note: 3G#Ab
	assign memory[	 51	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 52	] =	{1'd0, 6'd50, 6'd60, 3'd0};	// Note: 5A#Bb
	assign memory[	 53	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 54	] =	{1'd0, 6'd39, 6'd24, 3'd0};	// Note: 4B
	assign memory[	 55	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 56	] =	{1'd0, 6'd45, 6'd24, 3'd0};	// Note: 4F
	assign memory[	 57	] =	{1'd0, 6'd42, 6'd24, 3'd0};	// Note: 4D
	assign memory[	 58	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 59	] =	{1'd0, 6'd50, 6'd48, 3'd0};	// Note: 5A#Bb
	assign memory[	 60	] =	{1'd0, 6'd39, 6'd24, 3'd0};	// Note: 4B
	assign memory[	 61	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 62	] =	{1'd0, 6'd45, 6'd24, 3'd0};	// Note: 4F
	assign memory[	 63	] =	{1'd0, 6'd41, 6'd24, 3'd0};	// Note: 4C#Db
	assign memory[	 64	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 65	] =	{1'd0, 6'd33, 6'd24, 3'd0};	// Note: 3F
	assign memory[	 66	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 67	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	 68	] =	{1'd0, 6'd40, 6'd24, 3'd0};	// Note: 4C
	assign memory[	 69	] =	{1'd0, 6'd36, 6'd24, 3'd0};	// Note: 3G#Ab
	assign memory[	 70	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 71	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	 72	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 73	] =	{1'd0, 6'd48, 6'd12, 3'd0};	// Note: 4G#Ab
	assign memory[	 74	] =	{1'd0, 6'd33, 6'd24, 3'd0};	// Note: 3F
	assign memory[	 75	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 76	] =	{1'd0, 6'd48, 6'd12, 3'd0};	// Note: 4G#Ab
	assign memory[	 77	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 78	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	 79	] =	{1'd0, 6'd40, 6'd24, 3'd0};	// Note: 4C
	assign memory[	 80	] =	{1'd0, 6'd36, 6'd24, 3'd0};	// Note: 3G#Ab
	assign memory[	 81	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 82	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	 83	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 84	] =	{1'd0, 6'd52, 6'd12, 3'd0};	// Note: 5C
	assign memory[	 85	] =	{1'd0, 6'd36, 6'd24, 3'd0};	// Note: 3G#Ab
	assign memory[	 86	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 87	] =	{1'd0, 6'd52, 6'd24, 3'd0};	// Note: 5C
	assign memory[	 88	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 89	] =	{1'd0, 6'd43, 6'd24, 3'd0};	// Note: 4D#Eb
	assign memory[	 90	] =	{1'd0, 6'd40, 6'd24, 3'd0};	// Note: 4C
	assign memory[	 91	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 92	] =	{1'd0, 6'd52, 6'd24, 3'd0};	// Note: 5C
	assign memory[	 93	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 94	] =	{1'd0, 6'd36, 6'd24, 3'd0};	// Note: 3G#Ab
	assign memory[	 95	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 96	] =	{1'd0, 6'd48, 6'd12, 3'd0};	// Note: 4G#Ab
	assign memory[	 97	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	 98	] =	{1'd0, 6'd43, 6'd24, 3'd0};	// Note: 4D#Eb
	assign memory[	 99	] =	{1'd0, 6'd40, 6'd24, 3'd0};	// Note: 4C
	assign memory[	100	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	101	] =	{1'd0, 6'd50, 6'd12, 3'd0};	// Note: 5A#Bb
	assign memory[	102	] =	{1'd0, 6'd31, 6'd24, 3'd0};	// Note: 3D#Eb
	assign memory[	103	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	104	] =	{1'd0, 6'd50, 6'd24, 3'd0};	// Note: 5A#Bb
	assign memory[	105	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	106	] =	{1'd0, 6'd38, 6'd24, 3'd0};	// Note: 4A#Bb
	assign memory[	107	] =	{1'd0, 6'd35, 6'd24, 3'd0};	// Note: 3G
	assign memory[	108	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	109	] =	{1'd0, 6'd50, 6'd24, 3'd0};	// Note: 5A#Bb
	assign memory[	110	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	111	] =	{1'd0, 6'd31, 6'd24, 3'd0};	// Note: 3D#Eb
	assign memory[	112	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	113	] =	{1'd0, 6'd47, 6'd12, 3'd0};	// Note: 4G
	assign memory[	114	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	115	] =	{1'd0, 6'd38, 6'd24, 3'd0};	// Note: 4A#Bb
	assign memory[	116	] =	{1'd0, 6'd35, 6'd24, 3'd0};	// Note: 3G
	assign memory[	117	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	118	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	119	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	120	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	121	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	122	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	123	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	124	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	125	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	126	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	127	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	128	] =	{1'd0, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	129	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	130	] =	{1'd0, 6'd56, 6'd6, 3'd0};	// Note: 5E
	assign memory[	131	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	132	] =	{1'd0, 6'd54, 6'd6, 3'd0};	// Note: 5D#
	assign memory[	133	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	134	] =	{1'd0, 6'd56, 6'd6, 3'd0};	// Note: 5E
	assign memory[	135	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	136	] =	{1'd0, 6'd54, 6'd6, 3'd0};	// Note: 5D#
	assign memory[	137	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	138	] =	{1'd0, 6'd56, 6'd6, 3'd0};	// Note: 5E
	assign memory[	139	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	140	] =	{1'd0, 6'd51, 6'd6, 3'd0};	// Note: 5B
	assign memory[	141	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	142	] =	{1'd0, 6'd54, 6'd6, 3'd0};	// Note: 5D
	assign memory[	143	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	144	] =	{1'd0, 6'd52, 6'd6, 3'd0};	// Note: 5C
	assign memory[	145	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	146	] =	{1'd0, 6'd49, 6'd12, 3'd0};	// Note: 5A
	assign memory[	147	] =	{1'd0, 6'd37, 6'd24, 3'd0};	// Note: 4A
	assign memory[	148	] =	{1'd1, 6'd0, 6'd18, 3'd0};	// Note: rest
	assign memory[	149	] =	{1'd0, 6'd40, 6'd6, 3'd0};	// Note: 4C
	assign memory[	150	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	151	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	152	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	153	] =	{1'd0, 6'd49, 6'd6, 3'd0};	// Note: 5A
	assign memory[	154	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	155	] =	{1'd0, 6'd51, 6'd12, 3'd0};	// Note: 5B
	assign memory[	156	] =	{1'd0, 6'd32, 6'd24, 3'd0};	// Note: 3E
	assign memory[	157	] =	{1'd1, 6'd0, 6'd18, 3'd0};	// Note: rest
	assign memory[	158	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	159	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	160	] =	{1'd0, 6'd47, 6'd6, 3'd0};	// Note: 4G#
	assign memory[	161	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	162	] =	{1'd0, 6'd51, 6'd6, 3'd0};	// Note: 5B
	assign memory[	163	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	164	] =	{1'd0, 6'd52, 6'd12, 3'd0};	// Note: 5C
	assign memory[	165	] =	{1'd0, 6'd37, 6'd24, 3'd0};	// Note: 4A
	assign memory[	166	] =	{1'd1, 6'd0, 6'd18, 3'd0};	// Note: rest
	assign memory[	167	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	168	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	169	] =	{1'd0, 6'd56, 6'd6, 3'd0};	// Note: 5E
	assign memory[	170	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	171	] =	{1'd0, 6'd54, 6'd6, 3'd0};	// Note: 5D#
	assign memory[	172	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	173	] =	{1'd0, 6'd56, 6'd6, 3'd0};	// Note: 5E
	assign memory[	174	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	175	] =	{1'd0, 6'd54, 6'd6, 3'd0};	// Note: 5D#
	assign memory[	176	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	177	] =	{1'd0, 6'd56, 6'd6, 3'd0};	// Note: 5E
	assign memory[	178	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	179	] =	{1'd0, 6'd51, 6'd6, 3'd0};	// Note: 5B
	assign memory[	180	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	181	] =	{1'd0, 6'd54, 6'd6, 3'd0};	// Note: 5D
	assign memory[	182	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	183	] =	{1'd0, 6'd52, 6'd6, 3'd0};	// Note: 5C
	assign memory[	184	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	185	] =	{1'd0, 6'd49, 6'd12, 3'd0};	// Note: 5A
	assign memory[	186	] =	{1'd0, 6'd37, 6'd24, 3'd0};	// Note: 4A
	assign memory[	187	] =	{1'd1, 6'd0, 6'd18, 3'd0};	// Note: rest
	assign memory[	188	] =	{1'd0, 6'd40, 6'd6, 3'd0};	// Note: 4C
	assign memory[	189	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	190	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	191	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	192	] =	{1'd0, 6'd49, 6'd6, 3'd0};	// Note: 5A
	assign memory[	193	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	194	] =	{1'd0, 6'd51, 6'd12, 3'd0};	// Note: 5B
	assign memory[	195	] =	{1'd0, 6'd32, 6'd24, 3'd0};	// Note: 3E
	assign memory[	196	] =	{1'd1, 6'd0, 6'd18, 3'd0};	// Note: rest
	assign memory[	197	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	198	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	199	] =	{1'd0, 6'd52, 6'd6, 3'd0};	// Note: 5C
	assign memory[	200	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	201	] =	{1'd0, 6'd51, 6'd6, 3'd0};	// Note: 5B
	assign memory[	202	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	203	] =	{1'd0, 6'd49, 6'd12, 3'd0};	// Note: 5A
	assign memory[	204	] =	{1'd0, 6'd37, 6'd24, 3'd0};	// Note: 4A
	assign memory[	205	] =	{1'd1, 6'd0, 6'd18, 3'd0};	// Note: rest
	assign memory[	206	] =	{1'd0, 6'd51, 6'd6, 3'd0};	// Note: 5B
	assign memory[	207	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	208	] =	{1'd0, 6'd52, 6'd6, 3'd0};	// Note: 5C
	assign memory[	209	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	210	] =	{1'd0, 6'd54, 6'd6, 3'd0};	// Note: 5D
	assign memory[	211	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	212	] =	{1'd0, 6'd56, 6'd12, 3'd0};	// Note: 5E
	assign memory[	213	] =	{1'd0, 6'd40, 6'd24, 3'd0};	// Note: 4C
	assign memory[	214	] =	{1'd1, 6'd0, 6'd18, 3'd0};	// Note: rest
	assign memory[	215	] =	{1'd0, 6'd47, 6'd6, 3'd0};	// Note: 4G
	assign memory[	216	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	217	] =	{1'd0, 6'd57, 6'd6, 3'd0};	// Note: 5F
	assign memory[	218	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	219	] =	{1'd0, 6'd56, 6'd6, 3'd0};	// Note: 5E
	assign memory[	220	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	221	] =	{1'd0, 6'd54, 6'd12, 3'd0};	// Note: 5D
	assign memory[	222	] =	{1'd0, 6'd39, 6'd24, 3'd0};	// Note: 4B
	assign memory[	223	] =	{1'd1, 6'd0, 6'd18, 3'd0};	// Note: rest
	assign memory[	224	] =	{1'd0, 6'd45, 6'd6, 3'd0};	// Note: 4F
	assign memory[	225	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	226	] =	{1'd0, 6'd56, 6'd6, 3'd0};	// Note: 5E
	assign memory[	227	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	228	] =	{1'd0, 6'd54, 6'd6, 3'd0};	// Note: 5D
	assign memory[	229	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	230	] =	{1'd0, 6'd52, 6'd12, 3'd0};	// Note: 5C
	assign memory[	231	] =	{1'd0, 6'd37, 6'd24, 3'd0};	// Note: 4A
	assign memory[	232	] =	{1'd1, 6'd0, 6'd18, 3'd0};	// Note: rest
	assign memory[	233	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	234	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	235	] =	{1'd0, 6'd54, 6'd6, 3'd0};	// Note: 5D
	assign memory[	236	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	237	] =	{1'd0, 6'd52, 6'd6, 3'd0};	// Note: 5C
	assign memory[	238	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	239	] =	{1'd0, 6'd51, 6'd36, 3'd0};	// Note: 5B
	assign memory[	240	] =	{1'd0, 6'd35, 6'd36, 3'd0};	// Note: 3G#
	assign memory[	241	] =	{1'd1, 6'd0, 6'd36, 3'd0};	// Note: rest
	assign memory[	242	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	243	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	244	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	245	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	246	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	247	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	248	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	249	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	250	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	251	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	252	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	253	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	254	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	255	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	256	] =	{1'd0, 6'd47, 6'd48, 3'd0};	// Note: 4G
	assign memory[	257	] =	{1'd0, 6'd44, 6'd48, 3'd0};	// Note: 4E
	assign memory[	258	] =	{1'd0, 6'd40, 6'd48, 3'd0};	// Note: 4C
	assign memory[	259	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	260	] =	{1'd0, 6'd49, 6'd48, 3'd0};	// Note: 5A
	assign memory[	261	] =	{1'd0, 6'd45, 6'd48, 3'd0};	// Note: 4F
	assign memory[	262	] =	{1'd0, 6'd42, 6'd48, 3'd0};	// Note: 4D
	assign memory[	263	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	264	] =	{1'd0, 6'd51, 6'd48, 3'd0};	// Note: 5B
	assign memory[	265	] =	{1'd0, 6'd47, 6'd48, 3'd0};	// Note: 4G
	assign memory[	266	] =	{1'd0, 6'd44, 6'd48, 3'd0};	// Note: 4E
	assign memory[	267	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	268	] =	{1'd0, 6'd52, 6'd48, 3'd0};	// Note: 5C
	assign memory[	269	] =	{1'd0, 6'd49, 6'd48, 3'd0};	// Note: 5A
	assign memory[	270	] =	{1'd0, 6'd45, 6'd48, 3'd0};	// Note: 4F
	assign memory[	271	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	272	] =	{1'd0, 6'd54, 6'd48, 3'd0};	// Note: 5D
	assign memory[	273	] =	{1'd0, 6'd51, 6'd48, 3'd0};	// Note: 5B
	assign memory[	274	] =	{1'd0, 6'd47, 6'd48, 3'd0};	// Note: 4G
	assign memory[	275	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	276	] =	{1'd0, 6'd56, 6'd48, 3'd0};	// Note: 5E
	assign memory[	277	] =	{1'd0, 6'd52, 6'd48, 3'd0};	// Note: 5C
	assign memory[	278	] =	{1'd0, 6'd49, 6'd48, 3'd0};	// Note: 5A
	assign memory[	279	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	280	] =	{1'd0, 6'd57, 6'd48, 3'd0};	// Note: 5F
	assign memory[	281	] =	{1'd0, 6'd54, 6'd48, 3'd0};	// Note: 5D
	assign memory[	282	] =	{1'd0, 6'd51, 6'd48, 3'd0};	// Note: 5B
	assign memory[	283	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	284	] =	{1'd0, 6'd59, 6'd48, 3'd0};	// Note: 5G
	assign memory[	285	] =	{1'd0, 6'd56, 6'd48, 3'd0};	// Note: 5E
	assign memory[	286	] =	{1'd0, 6'd52, 6'd48, 3'd0};	// Note: 5C
	assign memory[	287	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	288	] =	{1'd0, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	289	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	290	] =	{1'd0, 6'd47, 6'd48, 3'd0};	// Note: 4G
	assign memory[	291	] =	{1'd0, 6'd43, 6'd48, 3'd0};	// Note: 4D#Eb
	assign memory[	292	] =	{1'd0, 6'd40, 6'd48, 3'd0};	// Note: 4C
	assign memory[	293	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	294	] =	{1'd0, 6'd48, 6'd48, 3'd0};	// Note: 4G#Ab
	assign memory[	295	] =	{1'd0, 6'd45, 6'd48, 3'd0};	// Note: 4F
	assign memory[	296	] =	{1'd0, 6'd42, 6'd48, 3'd0};	// Note: 4D
	assign memory[	297	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	298	] =	{1'd0, 6'd50, 6'd48, 3'd0};	// Note: 5A#Bb
	assign memory[	299	] =	{1'd0, 6'd47, 6'd48, 3'd0};	// Note: 4G
	assign memory[	300	] =	{1'd0, 6'd43, 6'd48, 3'd0};	// Note: 4D#Eb
	assign memory[	301	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	302	] =	{1'd0, 6'd52, 6'd48, 3'd0};	// Note: 5C
	assign memory[	303	] =	{1'd0, 6'd48, 6'd48, 3'd0};	// Note: 4G#Ab
	assign memory[	304	] =	{1'd0, 6'd45, 6'd48, 3'd0};	// Note: 4F
	assign memory[	305	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	306	] =	{1'd0, 6'd54, 6'd48, 3'd0};	// Note: 5D
	assign memory[	307	] =	{1'd0, 6'd50, 6'd48, 3'd0};	// Note: 5A#Bb
	assign memory[	308	] =	{1'd0, 6'd47, 6'd48, 3'd0};	// Note: 4G
	assign memory[	309	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	310	] =	{1'd0, 6'd55, 6'd48, 3'd0};	// Note: 5D#Eb
	assign memory[	311	] =	{1'd0, 6'd52, 6'd48, 3'd0};	// Note: 5C
	assign memory[	312	] =	{1'd0, 6'd48, 6'd48, 3'd0};	// Note: 4G#Ab
	assign memory[	313	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	314	] =	{1'd0, 6'd57, 6'd48, 3'd0};	// Note: 5F
	assign memory[	315	] =	{1'd0, 6'd54, 6'd48, 3'd0};	// Note: 5D
	assign memory[	316	] =	{1'd0, 6'd50, 6'd48, 3'd0};	// Note: 5A#Bb
	assign memory[	317	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	318	] =	{1'd0, 6'd59, 6'd48, 3'd0};	// Note: 5G
	assign memory[	319	] =	{1'd0, 6'd55, 6'd48, 3'd0};	// Note: 5D#Eb
	assign memory[	320	] =	{1'd0, 6'd52, 6'd48, 3'd0};	// Note: 5C
	assign memory[	321	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	322	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	323	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	324	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	325	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	326	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	327	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	328	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	329	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	330	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	331	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	332	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	333	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	334	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	335	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	336	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	337	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	338	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	339	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	340	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	341	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	342	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	343	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	344	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	345	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	346	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	347	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	348	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	349	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	350	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	351	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	352	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	353	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	354	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	355	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	356	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	357	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	358	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	359	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	360	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	361	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	362	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	363	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	364	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	365	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	366	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	367	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	368	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	369	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	370	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	371	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	372	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	373	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	374	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	375	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	376	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	377	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	378	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	379	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	380	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	381	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	382	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	383	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	384	] =	{1'd0, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	385	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	386	] =	{1'd0, 6'd44, 6'd12, 3'd0};	// Note: 4E
	assign memory[	387	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	388	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	389	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	390	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F#
	assign memory[	391	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	392	] =	{1'd0, 6'd47, 6'd6, 3'd0};	// Note: 4G
	assign memory[	393	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	394	] =	{1'd0, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	395	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	396	] =	{1'd0, 6'd47, 6'd6, 3'd0};	// Note: 4G
	assign memory[	397	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	398	] =	{1'd0, 6'd47, 6'd6, 3'd0};	// Note: 4G
	assign memory[	399	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	400	] =	{1'd0, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	401	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	402	] =	{1'd0, 6'd47, 6'd6, 3'd0};	// Note: 4G
	assign memory[	403	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	404	] =	{1'd0, 6'd47, 6'd6, 3'd0};	// Note: 4G
	assign memory[	405	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	406	] =	{1'd0, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	407	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	408	] =	{1'd0, 6'd49, 6'd12, 3'd0};	// Note: 5A
	assign memory[	409	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	410	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	411	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	412	] =	{1'd0, 6'd47, 6'd48, 3'd0};	// Note: 4G
	assign memory[	413	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	414	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	415	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	416	] =	{1'd0, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	417	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	418	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	419	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	420	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	421	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	422	] =	{1'd0, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	423	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	424	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	425	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	426	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	427	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	428	] =	{1'd0, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	429	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	430	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	431	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	432	] =	{1'd0, 6'd42, 6'd12, 3'd0};	// Note: 4D
	assign memory[	433	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	434	] =	{1'd0, 6'd44, 6'd60, 3'd0};	// Note: 4E
	assign memory[	435	] =	{1'd1, 6'd0, 6'd60, 3'd0};	// Note: rest
	assign memory[	436	] =	{1'd0, 6'd44, 6'd12, 3'd0};	// Note: 4E
	assign memory[	437	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	438	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	439	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	440	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F#
	assign memory[	441	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	442	] =	{1'd0, 6'd47, 6'd6, 3'd0};	// Note: 4G
	assign memory[	443	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	444	] =	{1'd0, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	445	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	446	] =	{1'd0, 6'd47, 6'd6, 3'd0};	// Note: 4G
	assign memory[	447	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	448	] =	{1'd0, 6'd47, 6'd6, 3'd0};	// Note: 4G
	assign memory[	449	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	450	] =	{1'd0, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	451	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	452	] =	{1'd0, 6'd47, 6'd6, 3'd0};	// Note: 4G
	assign memory[	453	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	454	] =	{1'd0, 6'd47, 6'd6, 3'd0};	// Note: 4G
	assign memory[	455	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	456	] =	{1'd0, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	457	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	458	] =	{1'd0, 6'd49, 6'd12, 3'd0};	// Note: 5A
	assign memory[	459	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	460	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	461	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	462	] =	{1'd0, 6'd47, 6'd48, 3'd0};	// Note: 4G
	assign memory[	463	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	464	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	465	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	466	] =	{1'd0, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	467	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	468	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	469	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	470	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	471	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	472	] =	{1'd0, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	473	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	474	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	475	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	476	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	477	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	478	] =	{1'd0, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	479	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	480	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	481	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	482	] =	{1'd0, 6'd42, 6'd12, 3'd0};	// Note: 4D
	assign memory[	483	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	484	] =	{1'd0, 6'd40, 6'd48, 3'd0};	// Note: 4C
	assign memory[	485	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
	assign memory[	486	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	487	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	488	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	489	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	490	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	491	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	492	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	493	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	494	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	495	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	496	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	497	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	498	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	499	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	500	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	501	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	502	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	503	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	504	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	505	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	506	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	507	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	508	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	509	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	510	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
	assign memory[	511	] =	{1'd1, 6'd0, 6'd0, 3'd0};	// Note: rest
endmodule					